`timescale 1ns / 1ps

module freq_div(
	clk_i,
	reset_i,	// sync high
	clk_o
	);
    
    input          clk_i;
	input          reset_i;
	output         clk_o;
    

endmodule
