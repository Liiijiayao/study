
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/11/08 11:25:42
// Design Name: 
// Module Name: freq_div_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module freq_div_tb();
 
	

	freq_div 
	freq_div (
		.clk_i					(), 
		.reset_i				(), 
		.clk_o					()
	);
endmodule